///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: Decoder_32
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////

module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Input: A (5-bit)
reg[4:0] A;
///////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////
// Output: Q (32-bit)
wire[31:0] Q;
///////////////////////////////////////////////////////////////////////////////////

Decoder_32 myDecoder(A, Q[0], Q[1], Q[2], Q[3], Q[4], Q[5], Q[6], Q[7], Q[8], Q[9], Q[10], Q[11], Q[12], Q[13], Q[14], Q[15], Q[16], Q[17], Q[18], Q[19], Q[20], Q[21], Q[22], Q[23], Q[24], Q[25], Q[26], Q[27], Q[28], Q[29], Q[30], Q[31]);

initial begin
////////////////////////////////////////////////////////////////////////
//  Testing: All 5-bit A values
for (A = 5'b00000; A <= 5'b11111; A = A + 5'b00001) begin
   $display("Testing: A=%b", A);
   #10;
   verifyEqual32(Q, 2**A);
   // You need this because the counter will reset to 0 otherwise
   if (A == 5'b11111) begin
    $display("All tests passed.");
    $stop;
   end
end
////////////////////////////////////////////////////////////////////////


end

endmodule